module fft_top(
	input clk
);

fft_butterfly fft_butterfly();

endmodule