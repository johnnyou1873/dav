module midiSong #(
	parameter BASE_SPEED = 50000000
)(
	input logic clk,
	input logic rst,
	input logic play,
	input logic en [0:4],
	output logic [7:0] out // 8-bit amplitude
);

	logic [19:0] freq [0:4];
	
	initial begin
		for (int i = 0; i < 5; i++) begin
			counter[i] <= 0;
		end
	end
	
	logic [11:0] counter [0:4];
	logic [7:0] tone [0:4];
	logic [31:0] millis;
	logic millisClk;
	
	// W = width of each tone[], OUTW = width of out[]
	localparam W    = 8;
	localparam OUTW = 8;

	// Compute full‐width sum and do some mixing
	wire [W+1:0] sum = 
		((en[0] ? tone[0]: '0) +
		(en[1] ? tone[1]: '0) +
		(en[2] ? (tone[2] >> 2) : '0) +
		(en[3] ? (tone[3] >> 2) : '0) +
		(en[4] ? (tone[4] >> 2) : '0));

	// sum/3 using (sum * 85) >> 8 (since 85/256 = 1/3 exactly for 8-bits)
	wire [W+1:0] avg = (sum * 85) >> 8;

	// if avg is bigger than max, clamp it
	assign out = (avg >= { {(OUTW){1'b1}} }) ?
								{ {(OUTW){1'b1}} } :
								avg[OUTW-1:0];

	sineGenerator #(.BASE_SPEED(BASE_SPEED)) voice0 (.clk(clk), .rst(rst), .freq(freq[0]), .out(tone[0]));
	sineGenerator #(.BASE_SPEED(BASE_SPEED)) voice1 (.clk(clk), .rst(rst), .freq(freq[1]), .out(tone[1]));
	sawtoothGenerator #(.BASE_SPEED(BASE_SPEED)) voice2 (.clk(clk), .rst(rst), .freq(freq[2]), .out(tone[2]));
	logic tone3_clk;
	clockDivider #(.BASE_SPEED(BASE_SPEED)) voice3 (.clk(clk), .rst(rst), .freq(freq[3]), .clk0(tone3_clk));
	assign tone[3] = tone3_clk ? 8'hFF : 8'h00;
	noiseGenerator #(.BASE_SPEED(BASE_SPEED)) voice4 (.clk(clk), .rst(rst), .freq(freq[4]), .out(tone[4]));
	clockDivider millisClock (.clk(clk), .rst(rst || ~play), .freq(1000), .clk0(millisClk)); // slow down millis due to framerate error
	
	always @(posedge millisClk or posedge rst or negedge play) begin
		if (rst || ~play) begin
			millis <= 0;
			for (int i = 0; i < 5; i++) begin
				counter[i] <= 0;
			end
		end else begin
			millis <= millis + 1; // purposefully overflow
			// Voice 0 (melody 1)
			if (counter[0] < $size(d1)-1 && millis == d1[counter[0]+1]) begin
				counter[0] <= counter[0] + 1;
			end
			// Voice 1 (melody 2)
			if (counter[1] < $size(d2)-1 && millis == d2[counter[1]+1]) begin
				counter[1] <= counter[1] + 1;
			end
			// Voice 2 (harmony 1)
			if (counter[2] < $size(d3)-1 && millis == d3[counter[2]+1]) begin
				counter[2] <= counter[2] + 1;
			end
			// Voice 3 (harmony 2)
			if (counter[3] < $size(d4)-1 && millis == d4[counter[3]+1]) begin
				counter[3] <= counter[3] + 1;
			end
			// Voice 4 (percussion)
			if (counter[4] < $size(d5)-1 && millis == d5[counter[4]+1]) begin
				counter[4] <= counter[4] + 1;
			end
		end
	end

	always_comb begin
		if (play) begin
			freq[0] = m1[counter[0]];
			freq[1] = m2[counter[1]];
			freq[2] = m3[counter[2]];
			freq[3] = m4[counter[3]];
			freq[4] = m5[counter[4]];
		end else begin
			for (int i = 0; i < 5; i++) begin
				freq[i] <= 0;
			end
		end
	end
	
	logic [31:0] d1[1310] = '{
		0,13913,14103,14130,14320,14347,14538,14565,14755,14782,15190,15217,15407,15434,15624,15652,16059,16086,16494,16521,16711,16739,16929,16956,17146,17173,17364,17391,17581,17608,17798,17826,18016,18043,18233,18260,18668,18695,18885,18913,19103,19130,19320,19347,19538,19565,19755,19782,19972,19999,20190,20217,20407,20434,20624,20652,20842,20869,21059,21086,21277,21304,21494,21521,21711,21739,22146,22173,22364,22391,22581,22608,23016,23043,23451,23478,23668,23695,23885,23913,24103,24130,24320,24347,24538,24565,24755,24782,24972,24999,25190,25217,25624,25652,25842,25869,26059,26086,26494,26521,26929,26956,27364,27391,27798,27826,28016,28043,28233,28260,28451,28478,28668,28695,29103,29130,29320,29347,29538,29565,29972,29999,30407,30434,30624,30652,30842,30869,31059,31086,31277,31304,31494,31521,31711,31739,31929,31956,32146,32173,32581,32608,32798,32826,33016,33043,33233,33260,33451,33478,33668,33695,33885,33912,34103,34130,34320,34347,34537,34565,34755,34782,34972,34999,35190,35217,35407,35434,35624,35652,36059,36086,36277,36304,36494,36521,36929,36956,37364,37391,37581,37608,37798,37826,38016,38043,38233,38260,38451,38478,38668,38695,38885,38912,39103,39130,39537,39565,39755,39782,39972,39999,40407,40434,40842,40869,41277,41304,41711,41739,41929,41956,42146,42173,42364,42391,42581,42608,43016,43043,43233,43260,43451,43478,43668,43695,43885,43912,44103,44130,44320,44347,44755,44782,44972,44999,45190,45217,45407,45434,45624,45652,45842,45869,46059,46086,46494,46521,46711,46739,46929,46956,47146,47173,47364,47391,47581,47608,47798,47826,48233,48260,48451,48478,48668,48695,48885,48912,49103,49130,49320,49347,49537,49565,49972,49999,50190,50217,50407,50434,50624,50652,50842,50869,51059,51086,51277,51304,51711,51739,51929,51956,52146,52173,52364,52391,52581,52608,52798,52826,53016,53043,53451,53478,53668,53695,53885,53912,54103,54130,54320,54347,54537,54565,54755,54782,55190,55217,55407,55434,55624,55652,55842,55869,56059,56086,56277,56304,56494,56521,56929,56956,57146,57173,57364,57391,57581,57608,57798,57826,58016,58043,58233,58260,58668,58695,58885,58912,59103,59130,59320,59347,59537,59565,59755,59782,59972,59999,60407,60434,60624,60652,60842,60869,61059,61086,61277,61304,61494,61521,61711,61739,62146,62173,62364,62391,62581,62608,62798,62825,63016,63043,63233,63260,63450,63478,63885,63912,64103,64130,64320,64347,64537,64565,64755,64782,64972,64999,65190,65217,65624,65652,65842,65869,66059,66086,66277,66304,66494,66521,66711,66739,66929,66956,67364,67391,67581,67608,67798,67825,68016,68043,68233,68260,68450,68478,68668,68695,68885,69130,69320,69347,69537,69565,69755,69782,69972,69999,70190,70217,70407,70434,70842,70869,71059,71086,71277,71304,71494,71521,71711,71739,71929,71956,72146,72173,72581,72608,72798,72825,73016,73043,73233,73260,73450,73478,73668,73695,73885,73912,74320,74347,74537,74565,74755,74782,74972,74999,75190,75217,75407,75434,75624,75652,76059,76086,76277,76304,76494,76521,76711,76739,76929,76956,77146,77173,77364,77391,77798,77825,78016,78043,78233,78260,78450,78478,78668,78695,78885,78912,79103,79130,79537,79565,79755,79782,79972,79999,80190,80217,80407,80434,80624,80652,80842,80869,81277,81304,81494,81521,81711,81739,81929,81956,82146,82173,82364,82391,82581,82608,83016,83043,83233,83260,83450,83478,83668,83695,83885,83912,84103,84130,84320,84347,84755,84782,84972,84999,85190,85217,85407,85434,85624,85652,85842,85869,86059,86086,86494,86521,86711,86739,86929,86956,87146,87173,87364,87391,87581,87608,87798,87825,88233,88260,88450,88478,88668,88695,88885,88912,89103,89130,89320,89347,89537,89565,89972,89999,90190,90217,90407,90434,90624,90652,90842,90869,91059,91086,91277,91304,91711,91739,91929,91956,92146,92173,92364,92391,92581,92608,92798,92825,93016,93043,93450,93478,93668,93695,93885,93912,94103,94130,94320,94347,94537,94565,94755,94782,95190,95217,95407,95434,95624,95652,95842,95869,96059,96086,96277,96304,96494,96521,96711,111299,111304,111489,111494,111521,111711,111738,111929,111956,112146,112173,112581,112608,112798,112825,113016,113043,113450,113478,113885,113912,114103,114130,114320,114347,114537,114565,114755,114782,114972,114999,115190,115217,115407,115434,115624,115652,116059,116086,116277,116304,116494,116521,116711,116738,116929,116956,117146,117173,117363,117391,117581,117608,117798,117825,118016,118043,118233,118260,118450,118478,118668,118695,118885,118912,119103,119130,119537,119565,119755,119782,119972,119999,120407,120434,120842,120869,121059,121086,121277,121304,121494,121521,121711,121738,121929,121956,122146,122173,122363,122391,122581,122608,123016,123043,123233,123260,123450,123478,123885,123912,124320,124347,124755,124782,125190,125217,125407,125434,125624,125651,125842,125869,126059,126086,126494,126521,126711,126738,126929,126956,127363,127391,127798,127825,128016,128043,128233,128260,128450,128478,128668,128695,128885,128912,129103,129130,129320,129347,129537,129565,129972,129999,130190,130217,130407,130434,130624,130651,130842,130869,131059,131086,131276,131304,131494,131521,131711,131738,131929,131956,132146,132173,132363,132391,132581,132608,132798,132825,133016,133043,133450,133478,133668,133695,133885,133912,134320,134347,134755,134782,134972,134999,135190,135217,135407,135434,135624,135651,135842,135869,136059,136086,136276,136304,136494,136521,136929,136956,137146,137173,137363,137391,137798,137825,138233,138260,138668,138695,139103,139130,139320,139347,139537,139565,139755,139782,139972,139999,140407,140434,140624,140651,140842,140869,141059,141086,141276,141304,141494,141521,141711,141738,142146,142173,142363,142391,142581,142608,142798,142825,143016,143043,143233,143260,143450,143478,143885,143912,144103,144130,144320,144347,144537,144565,144755,144782,144972,144999,145190,145217,145624,145651,145842,145869,146059,146086,146276,146304,146494,146521,146711,146738,146929,146956,147363,147391,147581,147608,147798,147825,148016,148043,148233,148260,148450,148478,148668,148695,149103,149130,149320,149347,149537,149565,149755,149782,149972,149999,150190,150217,150407,150434,150842,150869,151059,151086,151276,151304,151494,151521,151711,151738,151929,151956,152146,152173,152581,152608,152798,152825,153016,153043,153233,153260,153450,153478,153668,153695,153885,153912,154320,154347,154537,154565,154755,154782,154972,154999,155189,155217,155407,155434,155624,155651,156059,156086,156276,156304,156494,156521,156711,156738,156929,156956,157146,157173,157363,157391,157798,157825,158016,158043,158233,158260,158450,158478,158668,158695,158885,158912,159103,159130,159537,159564,159755,159782,159972,159999,160189,160217,160407,160434,160624,160651,160842,160869,161276,161304,161494,161521,161711,161738,161929,161956,162146,162173,162363,162391,162581,162608,163016,163043,163233,163260,163450,163478,163668,163695,163885,163912,164103,164130,164320,164347,164755,164782,164972,164999,165189,165217,165407,165434,165624,165651,165842,165869,166059,166086,166276,166521,166711,166738,166929,166956,167146,167173,167363,167391,167581,167608,167798,167825,168233,168260,168450,168478,168668,168695,168885,168912,169103,169130,169320,169347,169537,169564,169972,169999,170189,170217,170407,170434,170624,170651,170842,170869,171059,171086,171276,171304,171711,171738,171929,171956,172146,172173,172363,172391,172581,172608,172798,172825,173016,173043,173450,173478,173668,173695,173885,173912,174103,174130,174320,174347,174537,174564,174755,174782,175189,175217,175407,175434,175624,175651,175842,175869,176059,176086,176276,176304,176494,176521,176929,176956,177146,177173,177363,177391,177581,177608,177798,177825,178016,178043,178233,178260,178668,178695,178885,178912,179103,179130,179320,179347,179537,179564,179755,179782,179972,179999,180407,180434,180624,180651,180842,180869,181059,181086,181276,181304,181494,181521,181711,181738,182146,182173,182363,182391,182581,182608,182798,182825,183016,183043,183233,183260,183450,183478,183885,183912,184103,184130,184320,184347,184537,184564,184755,184782,184972,184999,185189,185217,185624,185651,185842,185869,186059,186086,186276,186304,186494,186521,186711,186738,186929,186956,187363,187391,187581,187608,187798,187825,188016,188043,188233,188260,188450,188477,188668,188695,189102,189130,189320,189347,189537,189564,189755,189782,189972,189999,190189,190217,190407,190434,190842,190869,191059,191086,191276,191304,191494,191521,191711,191738,191929,191956,192146,192173,192581,192608,192798,192825,193016,193043,193233,193260,193450,193477,193668,193695,193885,193912,194755,199999,199999,200004
	};
	
	logic [31:0] m1[1310] = '{
		0,311,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,349,0,311,0,293,0,349,0,311,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,369,0,415,0,466,0,311,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,349,0,311,0,293,0,349,0,311,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,369,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,466,0,554,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,466,0,554,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,622,0,698,0,739,0,698,0,622,0,554,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,466,0,554,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,466,0,554,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,622,0,698,0,739,0,698,0,622,0,554,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,311,311,0,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,349,0,311,0,293,0,349,0,311,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,369,0,415,0,466,0,311,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,349,0,311,0,293,0,349,0,311,0,349,0,369,0,415,0,466,0,622,0,554,0,466,0,311,0,466,0,415,0,369,0,349,0,311,0,349,0,369,0,415,0,466,0,415,0,369,0,349,0,369,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,466,0,554,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,466,0,554,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,277,0,311,0,349,0,369,0,415,0,466,0,311,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,415,0,466,0,554,0,622,0,466,0,415,0,466,0,622,0,698,0,739,0,698,0,622,0,554,0,466,0,415,0,466,0,415,0,369,0,349,0,277,0,311,0,415,0,466,0,587,0,659,0,493,0,440,0,493,0,440,0,493,0,587,0,659,0,493,0,440,0,493,0,440,0,493,0,440,0,391,0,369,0,293,0,329,0,293,0,329,0,369,0,391,0,440,0,493,0,329,0,440,0,493,0,587,0,659,0,493,0,440,0,493,0,440,0,493,0,587,0,659,0,493,0,440,0,493,0,440,0,493,0,440,0,391,0,369,0,293,0,329,0,293,0,329,0,369,0,391,0,440,0,493,0,329,0,440,0,493,0,587,0,659,0,493,0,440,0,493,0,440,0,493,0,587,0,659,0,493,0,440,0,493,0,440,0,493,0,440,0,391,0,369,0,293,0,329,0,293,0,329,0,369,0,391,0,440,0,493,0,329,0,440,0,493,0,587,0,659,0,493,0,440,0,493,0,440,0,493,0,587,0,659,0,493,0,440,0,493,0,659,0,739,0,783,0,739,0,659,0,587,0,493,0,440,0,493,0,440,0,391,0,369,0,293,0,329,0,0,0,0
	};
	
	logic [31:0] d2[1100] = '{
		0,27826,27989,28043,28206,28260,28423,28478,28641,28695,29076,29130,29293,29347,29510,29565,29945,29999,30380,30434,30597,30652,30815,30869,31032,31086,31249,31304,31467,31521,31684,31739,31902,31956,32119,32173,32554,32608,32771,32826,32989,33043,33206,33260,33423,33478,33641,33695,33858,33912,34076,34130,34293,34347,34510,34565,34728,34782,34945,34999,35162,35217,35380,35434,35597,35652,36032,36086,36249,36304,36467,36521,36902,36956,37336,37391,37554,37608,37771,37826,37989,38043,38206,38260,38423,38478,38641,38695,38858,38912,39076,39130,39510,39565,39728,39782,39945,39999,40380,40434,40815,40869,41249,41304,41684,41739,41902,41956,42119,42173,42336,42391,42554,42608,42989,43043,43206,43260,43423,43478,43641,43695,43858,43912,44076,44130,44293,44347,44728,44782,44945,44999,45162,45217,45380,45434,45597,45652,45815,45869,46032,46086,46467,46521,46684,46739,46902,46956,47119,47173,47336,47391,47554,47608,47771,47826,48206,48260,48423,48478,48641,48695,48858,48912,49076,49130,49293,49347,49510,49565,49945,49999,50162,50217,50380,50434,50597,50652,50815,50869,51032,51086,51249,51304,51684,51739,51902,51956,52119,52173,52336,52391,52554,52608,52771,52826,52989,53043,53423,53478,53641,53695,53858,53912,54076,54130,54293,54347,54510,54565,54728,54782,55162,55217,55380,55434,55597,55652,55815,55869,56032,56086,56249,56304,56467,56521,56902,56956,57119,57173,57336,57391,57554,57608,57771,57826,57989,58043,58206,58260,58641,58695,58858,58912,59076,59130,59293,59347,59510,59565,59728,59782,59945,59999,60380,60434,60597,60652,60815,60869,61032,61086,61249,61304,61467,61521,61684,61739,62119,62173,62336,62391,62554,62608,62771,62825,62989,63043,63206,63260,63423,63478,63858,63912,64075,64130,64293,64347,64510,64565,64728,64782,64945,64999,65162,65217,65597,65652,65815,65869,66032,66086,66249,66304,66467,66521,66684,66739,66902,66956,67336,67391,67554,67608,67771,67825,67989,68043,68206,68260,68423,68478,68641,68695,68858,69130,69293,69347,69510,69565,69728,69782,69945,69999,70162,70217,70380,70434,70815,70869,71032,71086,71249,71304,71467,71521,71684,71739,71902,71956,72119,72173,72554,72608,72771,72825,72989,73043,73206,73260,73423,73478,73641,73695,73858,73912,74293,74347,74510,74565,74728,74782,74945,74999,75162,75217,75380,75434,75597,75652,76032,76086,76249,76304,76467,76521,76684,76739,76902,76956,77119,77173,77336,77391,77771,77825,77989,78043,78206,78260,78423,78478,78641,78695,78858,78912,79075,79130,79510,79565,79728,79782,79945,79999,80162,80217,80380,80434,80597,80652,80815,80869,81249,81304,81467,81521,81684,81739,81902,81956,82119,82173,82336,82391,82554,82608,82989,83043,83206,83260,83423,83478,83641,83695,83858,83912,84075,84130,84293,84347,84728,84782,84945,84999,85162,85217,85380,85434,85597,85652,85815,85869,86032,86086,86467,86521,86684,86739,86902,86956,87119,87173,87336,87391,87554,87608,87771,87825,88206,88260,88423,88478,88641,88695,88858,88912,89075,89130,89293,89347,89510,89565,89945,89999,90162,90217,90380,90434,90597,90652,90815,90869,91032,91086,91249,91304,91684,91739,91902,91956,92119,92173,92336,92391,92554,92608,92771,92825,92988,93043,93423,93478,93641,93695,93858,93912,94075,94130,94293,94347,94510,94565,94728,94782,95162,95217,95380,95434,95597,95652,95815,95869,96032,96086,96249,96304,96467,96521,96684,125217,125380,125434,125597,125651,125815,125869,126032,126086,126467,126521,126684,126738,126901,126956,127336,127391,127771,127825,127988,128043,128206,128260,128423,128478,128641,128695,128858,128912,129075,129130,129293,129347,129510,129565,129945,129999,130162,130217,130380,130434,130597,130651,130815,130869,131032,131086,131249,131304,131467,131521,131684,131738,131901,131956,132119,132173,132336,132391,132554,132608,132771,132825,132988,133043,133423,133478,133641,133695,133858,133912,134293,134347,134728,134782,134945,134999,135162,135217,135380,135434,135597,135651,135815,135869,136032,136086,136249,136304,136467,136521,136901,136956,137119,137173,137336,137391,137771,137825,138206,138260,138641,138695,139075,139130,139293,139347,139510,139565,139728,139782,139945,139999,140380,140434,140597,140651,140815,140869,141032,141086,141249,141304,141467,141521,141684,141738,142119,142173,142336,142391,142554,142608,142771,142825,142988,143043,143206,143260,143423,143478,143858,143912,144075,144130,144293,144347,144510,144565,144728,144782,144945,144999,145162,145217,145597,145651,145815,145869,146032,146086,146249,146304,146467,146521,146684,146738,146901,146956,147336,147391,147554,147608,147771,147825,147988,148043,148206,148260,148423,148478,148641,148695,149075,149130,149293,149347,149510,149565,149728,149782,149945,149999,150162,150217,150380,150434,150815,150869,151032,151086,151249,151304,151467,151521,151684,151738,151901,151956,152119,152173,152554,152608,152771,152825,152988,153043,153206,153260,153423,153478,153641,153695,153858,153912,154293,154347,154510,154565,154728,154782,154945,154999,155162,155217,155380,155434,155597,155651,156032,156086,156249,156304,156467,156521,156684,156738,156901,156956,157119,157173,157336,157391,157771,157825,157988,158043,158206,158260,158423,158478,158641,158695,158858,158912,159075,159130,159510,159564,159728,159782,159945,159999,160162,160217,160380,160434,160597,160651,160814,160869,161249,161304,161467,161521,161684,161738,161901,161956,162119,162173,162336,162391,162554,162608,162988,163043,163206,163260,163423,163478,163641,163695,163858,163912,164075,164130,164293,164347,164728,164782,164945,164999,165162,165217,165380,165434,165597,165651,165814,165869,166032,166086,166467,166521,166684,166738,166901,166956,167119,167173,167336,167391,167554,167608,167771,167825,168206,168260,168423,168478,168641,168695,168858,168912,169075,169130,169293,169347,169510,169564,169945,169999,170162,170217,170380,170434,170597,170651,170814,170869,171032,171086,171249,171304,171684,171738,171901,171956,172119,172173,172336,172391,172554,172608,172771,172825,172988,173043,173423,173478,173641,173695,173858,173912,174075,174130,174293,174347,174510,174564,174728,174782,175162,175217,175380,175434,175597,175651,175814,175869,176032,176086,176249,176304,176467,176521,176901,176956,177119,177173,177336,177391,177554,177608,177771,177825,177988,178043,178206,178260,178641,178695,178858,178912,179075,179130,179293,179347,179510,179564,179728,179782,179945,179999,180380,180434,180597,180651,180814,180869,181032,181086,181249,181304,181467,181521,181684,181738,182119,182173,182336,182391,182554,182608,182771,182825,182988,183043,183206,183260,183423,183478,183858,183912,184075,184130,184293,184347,184510,184564,184728,184782,184945,184999,185162,185217,185597,185651,185814,185869,186032,186086,186249,186304,186467,186521,186684,186738,186901,186956,187336,187391,187554,187608,187771,187825,187988,188043,188206,188260,188423,188477,188641,188695,189075,189130,189293,189347,189510,189564,189727,189782,189945,189999,190162,190217,190380,190434,190814,190869,191032,191086,191249,191304,191467,191521,191684,191738,191901,191956,192119,192173,192554,192608,192771,192825,192988,193043,193206,193260,193423,193477,193641,193695,193858,193912,194727,199999,199999,200004
	};
	
	logic [31:0] m2[1100] = '{
		0,233,0,277,0,311,0,349,0,369,0,466,0,415,0,369,0,233,0,369,0,349,0,311,0,277,0,246,0,277,0,311,0,349,0,369,0,349,0,311,0,277,0,233,0,277,0,311,0,293,0,261,0,233,0,293,0,233,0,277,0,311,0,349,0,369,0,466,0,415,0,369,0,233,0,369,0,349,0,311,0,277,0,246,0,277,0,311,0,349,0,369,0,349,0,311,0,277,0,311,0,349,0,369,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,349,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,349,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,349,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,415,0,466,0,466,0,415,0,369,0,311,0,311,0,277,0,311,0,233,0,207,0,207,0,174,0,184,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,311,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,311,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,311,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,415,0,466,0,466,0,415,0,369,0,349,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,233,0,277,0,311,0,349,0,369,0,466,0,415,0,369,0,233,0,369,0,349,0,311,0,277,0,246,0,277,0,311,0,349,0,369,0,349,0,311,0,277,0,233,0,277,0,311,0,293,0,261,0,233,0,293,0,233,0,277,0,311,0,349,0,369,0,466,0,415,0,369,0,233,0,369,0,349,0,311,0,277,0,246,0,277,0,311,0,349,0,369,0,349,0,311,0,277,0,311,0,349,0,369,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,349,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,349,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,349,0,349,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,349,0,369,0,311,0,277,0,311,0,277,0,311,0,277,0,233,0,207,0,174,0,184,0,174,0,184,0,207,0,233,0,277,0,311,0,184,0,311,0,349,0,369,0,391,0,329,0,293,0,329,0,293,0,329,0,369,0,391,0,329,0,293,0,329,0,293,0,329,0,293,0,246,0,220,0,184,0,195,0,184,0,195,0,220,0,246,0,293,0,329,0,195,0,329,0,369,0,369,0,391,0,329,0,293,0,329,0,293,0,329,0,369,0,391,0,329,0,293,0,329,0,293,0,329,0,293,0,246,0,220,0,184,0,195,0,184,0,195,0,220,0,246,0,293,0,329,0,195,0,329,0,369,0,369,0,391,0,329,0,293,0,329,0,293,0,329,0,369,0,391,0,329,0,293,0,329,0,293,0,329,0,293,0,246,0,220,0,184,0,195,0,184,0,195,0,220,0,246,0,293,0,329,0,195,0,329,0,369,0,369,0,391,0,329,0,293,0,329,0,293,0,329,0,369,0,391,0,329,0,293,0,329,0,440,0,493,0,493,0,440,0,391,0,369,0,329,0,293,0,329,0,293,0,246,0,220,0,184,0,195,0,0,0,0
	};

	logic [31:0] d3[1902] = '{
		0,13913,14103,14130,14211,14239,14320,14456,14538,14565,14646,14673,14755,14782,14972,14999,15081,15108,15190,15326,15407,15434,15516,15543,15624,15652,15842,15869,15951,15978,16059,16195,16277,16304,16385,16413,16494,16521,16711,16739,16820,16847,16929,16956,17146,17173,17255,17282,17364,17391,17581,17608,17690,17717,17798,17934,18016,18043,18124,18152,18233,18260,18451,18478,18559,18586,18668,18804,18885,18913,18994,19021,19103,19130,19320,19347,19429,19456,19538,19673,19755,19782,19864,19891,19972,19999,20190,20217,20298,20326,20407,20434,20624,20652,20733,20760,20842,20869,21059,21086,21168,21195,21277,21413,21494,21521,21603,21630,21711,21739,21929,21956,22038,22065,22146,22282,22364,22391,22472,22499,22581,22608,22798,22826,22907,22934,23016,23152,23233,23260,23342,23369,23451,23478,23668,23695,23777,23804,23885,23913,24103,24130,24211,24239,24320,24347,24538,24565,24646,24673,24755,24891,24972,24999,25081,25108,25190,25217,25407,25434,25516,25543,25624,25760,25842,25869,25951,25978,26059,26086,26277,26304,26385,26413,26494,26630,26711,26739,26820,26847,26929,26956,27146,27173,27255,27282,27364,27391,27581,27608,27690,27717,27798,27826,28016,28043,28124,28152,28233,28369,28451,28478,28559,28586,28668,28695,28885,28913,28994,29021,29103,29239,29320,29347,29429,29456,29538,29565,29755,29782,29864,29891,29972,30108,30190,30217,30298,30326,30407,30434,30624,30652,30733,30760,30842,30869,31059,31086,31168,31195,31277,31304,31494,31521,31603,31630,31711,31847,31929,31956,32037,32065,32146,32173,32364,32391,32472,32499,32581,32717,32798,32826,32907,32934,33016,33043,33233,33260,33342,33369,33451,33586,33668,33695,33777,33804,33885,33912,34103,34130,34211,34239,34320,34347,34537,34565,34646,34673,34755,34782,34972,34999,35081,35108,35190,35326,35407,35434,35516,35543,35624,35652,35842,35869,35951,35978,36059,36195,36277,36304,36385,36412,36494,36521,36711,36739,36820,36847,36929,37065,37146,37173,37255,37282,37364,37391,37581,37608,37690,37717,37798,37826,38016,38043,38124,38152,38233,38260,38451,38478,38559,38586,38668,38804,38885,38912,38994,39021,39103,39130,39320,39347,39429,39456,39537,39673,39755,39782,39864,39891,39972,39999,40190,40217,40407,40434,40624,40652,40842,40869,41059,41086,41277,41304,41494,41521,41711,41739,41929,41956,42037,42065,42146,42282,42364,42391,42472,42499,42581,42608,42798,42826,42907,42934,43016,43152,43233,43260,43342,43369,43451,43478,43668,43695,43777,43804,43885,44021,44103,44130,44211,44239,44320,44347,44537,44565,44646,44673,44755,44891,44972,44999,45081,45108,45190,45217,45407,45434,45516,45543,45624,45760,45842,45869,45951,45978,46059,46086,46277,46304,46385,46412,46494,46630,46711,46739,46820,46847,46929,46956,47146,47173,47255,47282,47364,47499,47581,47608,47690,47717,47798,47826,48016,48043,48124,48152,48233,48260,48369,48451,48451,48478,48559,48586,48668,48695,48885,48912,48994,49021,49103,49239,49320,49347,49429,49456,49537,49565,49755,49782,49864,49891,49972,50108,50190,50217,50298,50326,50407,50434,50624,50652,50733,50760,50842,50978,51059,51086,51168,51195,51277,51304,51494,51521,51603,51630,51711,51847,51929,51956,52037,52065,52146,52173,52364,52391,52472,52499,52581,52717,52798,52826,52907,52934,53016,53043,53233,53260,53342,53369,53451,53586,53668,53695,53777,53804,53885,53912,54103,54130,54211,54239,54320,54456,54537,54565,54646,54673,54755,54782,54972,54999,55081,55108,55190,55217,55326,55407,55407,55434,55516,55543,55624,55652,55842,55869,55951,55978,56059,56195,56277,56304,56385,56412,56494,56521,56711,56739,56820,56847,56929,57065,57146,57173,57255,57282,57364,57391,57581,57608,57690,57717,57798,57934,58016,58043,58124,58152,58233,58260,58451,58478,58559,58586,58668,58804,58885,58912,58994,59021,59103,59130,59320,59347,59429,59456,59537,59673,59755,59782,59864,59891,59972,59999,60190,60217,60298,60326,60407,60543,60624,60652,60733,60760,60842,60869,61059,61086,61168,61195,61277,61412,61494,61521,61603,61630,61711,61739,61929,61956,62037,62065,62146,62173,62282,62364,62364,62391,62472,62499,62581,62608,62798,62825,62907,62934,63016,63152,63233,63260,63342,63369,63450,63478,63668,63695,63777,63804,63885,64021,64103,64130,64211,64239,64320,64347,64537,64565,64646,64673,64755,64891,64972,64999,65081,65108,65190,65217,65407,65434,65516,65543,65624,65760,65842,65869,65950,65978,66059,66086,66277,66304,66385,66412,66494,66630,66711,66739,66820,66847,66929,66956,67146,67173,67255,67282,67364,67499,67581,67608,67690,67717,67798,67825,68016,68043,68124,68152,68233,68369,68450,68478,68559,68586,68668,68695,68885,68912,68994,69021,69103,69130,69239,69320,69320,69347,69429,69456,69537,69565,71277,71304,73016,73043,76494,76521,78233,78260,79972,79999,83450,83478,85190,85217,86929,86956,90407,90434,92146,92173,93885,93912,95624,96521,96929,96956,97363,97391,97581,97608,97690,97717,97798,97934,98016,98043,98124,98152,98233,98260,98450,98478,98559,98586,98668,98804,98885,98912,98994,99021,99103,99130,99320,99347,99429,99456,99537,99673,99755,99782,99863,99891,99972,99999,100190,100217,100298,100325,100407,100434,100624,100652,100733,100760,100842,100869,101059,101086,101168,101195,101277,101412,101494,101521,101603,101630,101711,101738,101929,101956,102037,102065,102146,102282,102363,102391,102472,102499,102581,102608,102798,102825,102907,102934,103016,103152,103233,103260,103342,103369,103450,103478,103668,103695,103777,103804,103885,103912,104103,104130,104211,104238,104320,104347,104537,104565,104646,104673,104755,104891,104972,104999,105081,105108,105190,105217,105407,105434,105516,105543,105624,105760,105842,105869,105950,105978,106059,106086,106277,106304,106385,106412,106494,106630,106711,106738,106820,106847,106929,106956,107146,107173,107255,107282,107363,107391,107581,107608,107690,107717,107798,107825,108016,108043,108124,108152,108233,108369,108450,108478,108559,108586,108668,108695,108885,108912,108994,109021,109103,109238,109320,109347,109429,109456,109537,109565,109755,109782,109863,109891,109972,110108,110190,110217,110298,110325,110407,110434,110570,110597,110733,110760,110842,110869,111005,111005,111141,111168,111277,111304,111494,111521,111603,111630,111711,111847,111929,111956,112037,112065,112146,112173,112363,112391,112472,112499,112581,112717,112798,112825,112907,112934,113016,113043,113233,113260,113342,113369,113450,113586,113668,113695,113777,113804,113885,113912,114103,114130,114211,114238,114320,114347,114537,114565,114646,114673,114755,114782,114972,114999,115081,115108,115190,115325,115407,115434,115516,115543,115624,115652,115842,115869,115950,115978,116059,116195,116277,116304,116385,116412,116494,116521,116711,116738,116820,116847,116929,117065,117146,117173,117255,117282,117363,117391,117581,117608,117690,117717,117798,117825,118016,118043,118124,118152,118233,118260,118450,118478,118559,118586,118668,118804,118885,118912,118994,119021,119103,119130,119320,119347,119429,119456,119537,119673,119755,119782,119863,119891,119972,119999,120190,120217,120298,120325,120407,120543,120624,120652,120733,120760,120842,120869,121059,121086,121168,121195,121277,121304,121494,121521,121603,121630,121711,121738,121929,121956,122037,122065,122146,122282,122363,122391,122472,122499,122581,122608,122798,122825,122907,122934,123016,123152,123233,123260,123342,123369,123450,123478,123668,123695,123777,123804,123885,124021,124103,124130,124211,124238,124320,124347,124537,124565,124646,124673,124755,124782,124972,124999,125081,125108,125190,125217,125407,125434,125516,125543,125624,125760,125842,125869,125950,125978,126059,126086,126276,126304,126385,126412,126494,126630,126711,126738,126820,126847,126929,126956,127146,127173,127255,127282,127363,127499,127581,127608,127690,127717,127798,127825,128016,128043,128124,128151,128233,128260,128450,128478,128559,128586,128668,128695,128885,128912,128994,129021,129103,129238,129320,129347,129429,129456,129537,129565,129755,129782,129863,129891,129972,130108,130190,130217,130298,130325,130407,130434,130624,130651,130733,130760,130842,130978,131059,131086,131168,131195,131276,131304,131494,131521,131603,131630,131711,131738,131929,131956,132037,132065,132146,132173,132363,132391,132472,132499,132581,132717,132798,132825,132907,132934,133016,133043,133233,133260,133342,133369,133450,133586,133668,133695,133776,133804,133885,133912,134103,134130,134211,134238,134320,134456,134537,134565,134646,134673,134755,134782,134972,134999,135081,135108,135190,135217,135407,135434,135516,135543,135624,135651,135842,135869,135950,135978,136059,136195,136276,136304,136385,136412,136494,136521,136711,136738,136820,136847,136929,137065,137146,137173,137255,137282,137363,137391,137581,137608,137690,137717,137798,137934,138016,138043,138124,138151,138233,138260,138450,138478,138559,138586,138668,138695,138885,138912,138994,139021,139103,139130,139320,139347,139429,139456,139537,139673,139755,139782,139863,139891,139972,139999,140190,140217,140298,140325,140407,140543,140624,140651,140733,140760,140842,140869,141059,141086,141168,141195,141276,141412,141494,141521,141603,141630,141711,141738,141929,141956,142037,142065,142146,142282,142363,142391,142472,142499,142581,142608,142798,142825,142907,142934,143016,143151,143233,143260,143342,143369,143450,143478,143668,143695,143776,143804,143885,144021,144103,144130,144211,144238,144320,144347,144537,144565,144646,144673,144755,144891,144972,144999,145081,145108,145190,145217,145407,145434,145516,145543,145624,145651,145760,145842,145842,145869,145950,145978,146059,146086,146276,146304,146385,146412,146494,146630,146711,146738,146820,146847,146929,146956,147146,147173,147255,147282,147363,147499,147581,147608,147690,147717,147798,147825,148016,148043,148124,148151,148233,148369,148450,148478,148559,148586,148668,148695,148885,148912,148994,149021,149103,149238,149320,149347,149429,149456,149537,149565,149755,149782,149863,149891,149972,150108,150190,150217,150298,150325,150407,150434,150624,150651,150733,150760,150842,150978,151059,151086,151168,151195,151276,151304,151494,151521,151603,151630,151711,151847,151929,151956,152037,152065,152146,152173,152363,152391,152472,152499,152581,152608,152717,152798,152798,152825,152907,152934,153016,153043,153233,153260,153342,153369,153450,153586,153668,153695,153776,153804,153885,153912,154103,154130,154211,154238,154320,154456,154537,154565,154646,154673,154755,154782,154972,154999,155081,155108,155189,155325,155407,155434,155516,155543,155624,155651,155842,155869,155950,155978,156059,156195,156276,156304,156385,156412,156494,156521,156711,156738,156820,156847,156929,157064,157146,157173,157255,157282,157363,157391,157581,157608,157689,157717,157798,157934,158016,158043,158124,158151,158233,158260,158450,158478,158559,158586,158668,158804,158885,158912,158994,159021,159103,159130,159320,159347,159429,159456,159537,159564,159673,159755,159755,159782,159863,159891,159972,159999,160189,160217,160298,160325,160407,160543,160624,160651,160733,160760,160842,160869,161059,161086,161168,161195,161276,161412,161494,161521,161603,161630,161711,161738,161929,161956,162037,162064,162146,162282,162363,162391,162472,162499,162581,162608,162798,162825,162907,162934,163016,163151,163233,163260,163342,163369,163450,163478,163668,163695,163776,163804,163885,164021,164103,164130,164211,164238,164320,164347,164537,164564,164646,164673,164755,164891,164972,164999,165081,165108,165189,165217,165407,165434,165516,165543,165624,165760,165842,165869,165950,165978,166059,166086,166276,166304,166385,166412,166494,166521,166630,166711,166711,166738,166820,166847,166929,166956,168668,168695,170407,170434,173885,173912,175624,175651,177363,177391,180842,180869,181059,181086,181385,181412,181711,181738,181929,181956,182255,182282,182581,182608,182798,182825,183124,183151,183450,183478,183668,183695,183994,184021,184320,184347,184537,184564,184863,184891,185189,185217,185407,185434,185733,185760,186059,186086,186276,186304,186603,186630,186929,186956,187146,187173,187472,187499,187798,187825,188016,188043,188342,188369,188668,188695,188885,188912,189211,189238,189537,189564,189755,189782,190081,190108,190407,190434,190624,190651,190950,190977,191276,191304,191494,191521,191820,191847,192146,192173,192363,192391,192689,192717,193016,193043,193233,193260,193559,193586,193885,193912,194102,194130,194429,194456,194755,194782,194972,194999,195298,195325,195624,195651,195842,195869,196168,196195,196494,196521,196711,196738,197037,197064,197363,197391,197581,197608,197907,197934,198233,198260,198559,199999,199999,200004
	};

	logic [31:0] m3[1902] = '{
		0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,138,0,77,0,155,0,87,0,174,0,92,0,184,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,92,0,103,0,116,0,92,0,103,0,116,0,92,0,103,0,116,0,92,0,103,0,116,0,207,0,184,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,61,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,69,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,77,0,155,0,155,0,155,0,138,0,155,0,103,0,155,0,155,0,92,155,0,0,138,0,155,0,97,0,110,0,123,0,97,0,110,0,123,0,97,0,97,0,97,0,97,0,97,0,97,0,110,0,110,0,110,0,110,0,110,0,110,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,97,0,97,0,97,0,97,0,97,0,97,0,110,0,110,0,110,0,110,0,110,0,110,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,110,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,123,0,0,0,0
	};

	logic [31:0] d4[2085] = '{
		0,190,217,298,326,407,543,624,652,733,760,842,869,1059,1086,1168,1195,1277,1413,1494,1521,1603,1630,1711,1739,1929,1956,2038,2065,2146,2282,2364,2391,2472,2499,2581,2608,2798,2826,2907,2934,3016,3043,3233,3260,3342,3369,3451,3478,3668,3695,3777,3804,3885,4021,4103,4130,4211,4239,4320,4347,4538,4565,4646,4673,4755,4891,4972,4999,5081,5108,5190,5217,5407,5434,5516,5543,5624,5760,5842,5869,5951,5978,6059,6086,6277,6304,6385,6413,6494,6521,6711,6739,6820,6847,6929,6956,7146,7173,7255,7282,7364,7499,7581,7608,7690,7717,7798,7826,8016,8043,8124,8152,8233,8369,8451,8478,8559,8586,8668,8695,8885,8913,8994,9021,9103,9239,9320,9347,9429,9456,9538,9565,9755,9782,9864,9891,9972,9999,10190,10217,10298,10326,10407,10434,10624,10652,10733,10760,10842,10978,11059,11086,11168,11195,11277,11304,11494,11521,11603,11630,11711,11847,11929,11956,12038,12065,12146,12173,12364,12391,12472,12499,12581,12717,12798,12826,12907,12934,13016,13043,13233,13260,13342,13369,13451,13478,13668,13695,13777,13804,13885,13913,14103,14130,14211,14239,14320,14456,14538,14565,14646,14673,14755,14782,14972,14999,15081,15108,15190,15326,15407,15434,15516,15543,15624,15652,15842,15869,15951,15978,16059,16195,16277,16304,16385,16413,16494,16521,16711,16739,16820,16847,16929,16956,17146,17173,17255,17282,17364,17391,17581,17608,17690,17717,17798,17934,18016,18043,18124,18152,18233,18260,18451,18478,18559,18586,18668,18804,18885,18913,18994,19021,19103,19130,19320,19347,19429,19456,19538,19673,19755,19782,19864,19891,19972,19999,20190,20217,20298,20326,20407,20543,20624,20652,20733,20760,20842,20869,21059,21086,21168,21195,21277,21413,21494,21521,21603,21630,21711,21739,21929,21956,22038,22065,22146,22282,22364,22391,22472,22499,22581,22608,22798,22826,22907,22934,23016,23152,23233,23260,23342,23369,23451,23478,23668,23695,23777,23804,23885,23913,24103,24130,24211,24239,24320,24347,24538,24565,24646,24673,24755,24891,24972,24999,25081,25108,25190,25217,25407,25434,25516,25543,25624,25760,25842,25869,25951,25978,26059,26086,26277,26304,26385,26413,26494,26630,26711,26739,26820,26847,26929,26956,27146,27173,27255,27282,27364,27499,27581,27608,27690,27717,27798,27826,28016,28043,28124,28152,28233,28369,28451,28478,28559,28586,28668,28695,28885,28913,28994,29021,29103,29239,29320,29347,29429,29456,29538,29565,29755,29782,29864,29891,29972,30108,30190,30217,30298,30326,30407,30434,30624,30652,30733,30760,30842,30869,31059,31086,31168,31195,31277,31304,31494,31521,31603,31630,31711,31847,31929,31956,32037,32065,32146,32173,32364,32391,32472,32499,32581,32717,32798,32826,32907,32934,33016,33043,33233,33260,33342,33369,33451,33586,33668,33695,33777,33804,33885,33912,34103,34130,34211,34239,34320,34456,34537,34565,34646,34673,34755,34782,34972,34999,35081,35108,35190,35326,35407,35434,35516,35543,35624,35652,35842,35869,35951,35978,36059,36195,36277,36304,36385,36412,36494,36521,36711,36739,36820,36847,36929,37065,37146,37173,37255,37282,37364,37391,37581,37608,37690,37717,37798,37826,38016,38043,38124,38152,38233,38260,38451,38478,38559,38586,38668,38804,38885,38912,38994,39021,39103,39130,39320,39347,39429,39456,39537,39673,39755,39782,39864,39891,39972,39999,40190,40217,40298,40326,40407,40543,40624,40652,40733,40760,40842,40869,41059,41086,41168,41195,41277,41412,41494,41521,41603,41630,41711,41739,41929,41956,42037,42065,42146,42282,42364,42391,42472,42499,42581,42608,42798,42826,42907,42934,43016,43152,43233,43260,43342,43369,43451,43478,43668,43695,43777,43804,43885,44021,44103,44130,44211,44239,44320,44347,44537,44565,44646,44673,44755,44891,44972,44999,45081,45108,45190,45217,45407,45434,45516,45543,45624,45760,45842,45869,45951,45978,46059,46086,46277,46304,46385,46412,46494,46630,46711,46739,46820,46847,46929,46956,47146,47173,47255,47282,47364,47499,47581,47608,47690,47717,47798,47826,48016,48043,48124,48152,48233,48260,48451,48478,48559,48586,48668,48695,48885,48912,48994,49021,49103,49239,49320,49347,49429,49456,49537,49565,49755,49782,49864,49891,49972,50108,50190,50217,50298,50326,50407,50434,50624,50652,50733,50760,50842,50978,51059,51086,51168,51195,51277,51304,51494,51521,51603,51630,51711,51847,51929,51956,52037,52065,52146,52173,52364,52391,52472,52499,52581,52717,52798,52826,52907,52934,53016,53043,53233,53260,53342,53369,53451,53586,53668,53695,53777,53804,53885,53912,54103,54130,54211,54239,54320,54456,54537,54565,54646,54673,54755,54782,54972,54999,55081,55108,55190,55217,55407,55434,55516,55543,55624,55652,55842,55869,55951,55978,56059,56195,56277,56304,56385,56412,56494,56521,56711,56739,56820,56847,56929,57065,57146,57173,57255,57282,57364,57391,57581,57608,57690,57717,57798,57934,58016,58043,58124,58152,58233,58260,58451,58478,58559,58586,58668,58804,58885,58912,58994,59021,59103,59130,59320,59347,59429,59456,59537,59673,59755,59782,59864,59891,59972,59999,60190,60217,60298,60326,60407,60543,60624,60652,60733,60760,60842,60869,61059,61086,61168,61195,61277,61412,61494,61521,61603,61630,61711,61739,61929,61956,62037,62065,62146,62173,62364,62391,62472,62499,62581,62608,62798,62825,62907,62934,63016,63152,63233,63260,63342,63369,63450,63478,63668,63695,63777,63804,63885,64021,64103,64130,64211,64239,64320,64347,64537,64565,64646,64673,64755,64891,64972,64999,65081,65108,65190,65217,65407,65434,65516,65543,65624,65760,65842,65869,65950,65978,66059,66086,66277,66304,66385,66412,66494,66630,66711,66739,66820,66847,66929,66956,67146,67173,67255,67282,67364,67499,67581,67608,67690,67717,67798,67825,68016,68043,68124,68152,68233,68369,68450,68478,68559,68586,68668,68695,68885,68912,68994,69021,69103,69130,69320,69347,69429,69456,69537,69565,71277,71304,73016,73043,76494,76521,78233,78260,79972,79999,83450,83478,85190,85217,86929,86956,90407,90434,92146,92173,93885,93912,95624,96521,96929,96956,97363,97391,97581,97608,97690,97717,97798,97934,98016,98043,98124,98152,98233,98260,98450,98478,98559,98586,98668,98804,98885,98912,98994,99021,99103,99130,99320,99347,99429,99456,99537,99673,99755,99782,99863,99891,99972,99999,100190,100217,100298,100325,100407,100434,100624,100652,100733,100760,100842,100869,101059,101086,101168,101195,101277,101412,101494,101521,101603,101630,101711,101738,101929,101956,102037,102065,102146,102282,102363,102391,102472,102499,102581,102608,102798,102825,102907,102934,103016,103152,103233,103260,103342,103369,103450,103478,103668,103695,103777,103804,103885,103912,104103,104130,104211,104238,104320,104347,104537,104565,104646,104673,104755,104891,104972,104999,105081,105108,105190,105217,105407,105434,105516,105543,105624,105760,105842,105869,105950,105978,106059,106086,106277,106304,106385,106412,106494,106630,106711,106738,106820,106847,106929,106956,107146,107173,107255,107282,107363,107391,107581,107608,107690,107717,107798,107825,108016,108043,108124,108152,108233,108369,108450,108478,108559,108586,108668,108695,108885,108912,108994,109021,109103,109238,109320,109347,109429,109456,109537,109565,109755,109782,109863,109891,109972,110108,110190,110217,110298,110325,110407,110434,110570,110597,110733,110760,110842,110869,111005,111032,111168,111168,111277,111304,111494,111521,111603,111630,111711,111847,111929,111956,112037,112065,112146,112173,112363,112391,112472,112499,112581,112717,112798,112825,112907,112934,113016,113043,113233,113260,113342,113369,113450,113586,113668,113695,113777,113804,113885,113912,114103,114130,114211,114238,114320,114347,114537,114565,114646,114673,114755,114782,114972,114999,115081,115108,115190,115325,115407,115434,115516,115543,115624,115652,115842,115869,115950,115978,116059,116195,116277,116304,116385,116412,116494,116521,116711,116738,116820,116847,116929,117065,117146,117173,117255,117282,117363,117391,117581,117608,117690,117717,117798,117934,118016,118043,118124,118152,118233,118260,118450,118478,118559,118586,118668,118804,118885,118912,118994,119021,119103,119130,119320,119347,119429,119456,119537,119673,119755,119782,119863,119891,119972,119999,120190,120217,120298,120325,120407,120543,120624,120652,120733,120760,120842,120869,121059,121086,121168,121195,121277,121304,121494,121521,121603,121630,121711,121738,121929,121956,122037,122065,122146,122282,122363,122391,122472,122499,122581,122608,122798,122825,122907,122934,123016,123152,123233,123260,123342,123369,123450,123478,123668,123695,123777,123804,123885,124021,124103,124130,124211,124238,124320,124347,124537,124565,124646,124673,124755,124891,124972,124999,125081,125108,125190,125217,125407,125434,125516,125543,125624,125760,125842,125869,125950,125978,126059,126086,126276,126304,126385,126412,126494,126630,126711,126738,126820,126847,126929,126956,127146,127173,127255,127282,127363,127499,127581,127608,127690,127717,127798,127825,128016,128043,128124,128151,128233,128260,128450,128478,128559,128586,128668,128695,128885,128912,128994,129021,129103,129238,129320,129347,129429,129456,129537,129565,129755,129782,129863,129891,129972,130108,130190,130217,130298,130325,130407,130434,130624,130651,130733,130760,130842,130978,131059,131086,131168,131195,131276,131304,131494,131521,131603,131630,131711,131847,131929,131956,132037,132065,132146,132173,132363,132391,132472,132499,132581,132717,132798,132825,132907,132934,133016,133043,133233,133260,133342,133369,133450,133586,133668,133695,133776,133804,133885,133912,134103,134130,134211,134238,134320,134456,134537,134565,134646,134673,134755,134782,134972,134999,135081,135108,135190,135217,135407,135434,135516,135543,135624,135651,135842,135869,135950,135978,136059,136195,136276,136304,136385,136412,136494,136521,136711,136738,136820,136847,136929,137065,137146,137173,137255,137282,137363,137391,137581,137608,137690,137717,137798,137934,138016,138043,138124,138151,138233,138260,138450,138478,138559,138586,138668,138804,138885,138912,138994,139021,139103,139130,139320,139347,139429,139456,139537,139673,139755,139782,139863,139891,139972,139999,140190,140217,140298,140325,140407,140543,140624,140651,140733,140760,140842,140869,141059,141086,141168,141195,141276,141412,141494,141521,141603,141630,141711,141738,141929,141956,142037,142065,142146,142282,142363,142391,142472,142499,142581,142608,142798,142825,142907,142934,143016,143151,143233,143260,143342,143369,143450,143478,143668,143695,143776,143804,143885,144021,144103,144130,144211,144238,144320,144347,144537,144565,144646,144673,144755,144891,144972,144999,145081,145108,145190,145217,145407,145434,145516,145543,145624,145651,145842,145869,145950,145978,146059,146086,146276,146304,146385,146412,146494,146630,146711,146738,146820,146847,146929,146956,147146,147173,147255,147282,147363,147499,147581,147608,147690,147717,147798,147825,148016,148043,148124,148151,148233,148369,148450,148478,148559,148586,148668,148695,148885,148912,148994,149021,149103,149238,149320,149347,149429,149456,149537,149565,149755,149782,149863,149891,149972,150108,150190,150217,150298,150325,150407,150434,150624,150651,150733,150760,150842,150978,151059,151086,151168,151195,151276,151304,151494,151521,151603,151630,151711,151847,151929,151956,152037,152065,152146,152173,152363,152391,152472,152499,152581,152608,152798,152825,152907,152934,153016,153043,153233,153260,153342,153369,153450,153586,153668,153695,153776,153804,153885,153912,154103,154130,154211,154238,154320,154456,154537,154565,154646,154673,154755,154782,154972,154999,155081,155108,155189,155325,155407,155434,155516,155543,155624,155651,155842,155869,155950,155978,156059,156195,156276,156304,156385,156412,156494,156521,156711,156738,156820,156847,156929,157064,157146,157173,157255,157282,157363,157391,157581,157608,157689,157717,157798,157934,158016,158043,158124,158151,158233,158260,158450,158478,158559,158586,158668,158804,158885,158912,158994,159021,159103,159130,159320,159347,159429,159456,159537,159564,159755,159782,159863,159891,159972,159999,160189,160217,160298,160325,160407,160543,160624,160651,160733,160760,160842,160869,161059,161086,161168,161195,161276,161412,161494,161521,161603,161630,161711,161738,161929,161956,162037,162064,162146,162282,162363,162391,162472,162499,162581,162608,162798,162825,162907,162934,163016,163151,163233,163260,163342,163369,163450,163478,163668,163695,163776,163804,163885,164021,164103,164130,164211,164238,164320,164347,164537,164564,164646,164673,164755,164891,164972,164999,165081,165108,165189,165217,165407,165434,165516,165543,165624,165760,165842,165869,165950,165978,166059,166086,166276,166304,166385,166412,166494,166521,166711,166738,166820,166847,166929,166956,168668,168695,170407,170434,173885,173912,175624,175651,177363,177391,180842,180869,181059,181086,181385,181412,181711,181738,181929,181956,182255,182282,182581,182608,182798,182825,183124,183151,183450,183478,183668,183695,183994,184021,184320,184347,184537,184564,184863,184891,185189,185217,185407,185434,185733,185760,186059,186086,186276,186304,186603,186630,186929,186956,187146,187173,187472,187499,187798,187825,188016,188043,188342,188369,188668,188695,188885,188912,189211,189238,189537,189564,189755,189782,190081,190108,190407,190434,190624,190651,190950,190977,191276,191304,191494,191521,191820,191847,192146,192173,192363,192391,192689,192717,193016,193043,193233,193260,193559,193586,193885,193912,194102,194130,194429,194456,194755,194782,194972,194999,195298,195325,195624,195651,195842,195869,196168,196195,196494,196521,196711,196738,197037,197064,197363,197391,197581,197608,197907,197934,198233,198260,198559,199999,199999,200004
	};

	logic [31:0] m4[2085] = '{
		77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,61,0,69,0,77,0,61,0,69,0,77,0,61,0,69,0,77,0,61,0,69,0,77,0,103,0,92,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,155,0,184,0,103,0,184,0,207,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,73,0,73,0,146,0,146,0,116,0,146,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,61,0,61,0,123,0,123,0,116,0,123,0,61,0,61,0,123,0,123,0,116,0,123,0,69,0,69,0,138,0,138,0,123,0,138,0,69,0,69,0,138,0,138,0,123,0,138,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,77,0,77,0,155,0,155,0,138,0,155,0,103,0,184,0,207,0,92,0,155,0,184,0,65,0,73,0,82,0,65,0,73,0,82,0,65,0,65,0,65,0,65,0,65,0,65,0,73,0,73,0,73,0,73,0,73,0,73,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,65,0,65,0,65,0,65,0,65,0,65,0,73,0,73,0,73,0,73,0,73,0,73,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,73,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,82,0,0,0,0
	};

	logic [31:0] d5[1880] = '{
		0,6956,7146,7173,7255,7282,7364,7499,7581,7608,7690,7717,7798,7826,8016,8043,8124,8152,8233,8369,8451,8478,8559,8586,8668,8695,8885,8913,8994,9021,9103,9239,9320,9347,9429,9456,9538,9565,9755,9782,9864,9891,9972,9999,10190,10217,10298,10326,10407,10434,10624,10652,10733,10760,10842,10978,11059,11086,11168,11195,11277,11304,11494,11521,11603,11630,11711,11847,11929,11956,12038,12065,12146,12173,12364,12391,12472,12499,12581,12717,12798,12826,12907,12934,13016,13043,13233,13260,13342,13369,13451,13478,13668,13695,13777,13804,13885,13913,14103,14130,14211,14239,14320,14456,14538,14565,14646,14673,14755,14782,14972,14999,15081,15108,15190,15326,15407,15434,15516,15543,15624,15652,15842,15869,15951,15978,16059,16195,16277,16304,16385,16413,16494,16521,16711,16739,16820,16847,16929,16956,17146,17173,17255,17282,17364,17391,17581,17608,17690,17717,17798,17934,18016,18043,18124,18152,18233,18260,18451,18478,18559,18586,18668,18804,18885,18913,18994,19021,19103,19130,19320,19347,19429,19456,19538,19673,19755,19782,19864,19891,19972,19999,20190,20217,20298,20326,20407,20543,20624,20652,20733,20760,20842,20869,21059,21086,21168,21195,21277,21413,21494,21521,21603,21630,21711,21739,21929,21956,22038,22065,22146,22282,22364,22391,22472,22499,22581,22608,22798,22826,22907,22934,23016,23152,23233,23260,23342,23369,23451,23478,23668,23695,23777,23804,23885,23913,24103,24130,24211,24239,24320,24347,24538,24565,24646,24673,24755,24891,24972,24999,25081,25108,25190,25217,25407,25434,25516,25543,25624,25760,25842,25869,25951,25978,26059,26086,26277,26304,26385,26413,26494,26630,26711,26739,26820,26847,26929,26956,27146,27173,27255,27282,27364,27499,27581,27608,27690,27717,27798,27826,28016,28043,28124,28152,28233,28369,28451,28478,28559,28586,28668,28695,28885,28913,28994,29021,29103,29239,29320,29347,29429,29456,29538,29565,29755,29782,29864,29891,29972,30108,30190,30217,30298,30326,30407,30434,30624,30652,30733,30760,30842,30869,31059,31086,31168,31195,31277,31304,31494,31521,31603,31630,31711,31847,31929,31956,32037,32065,32146,32173,32364,32391,32472,32499,32581,32717,32798,32826,32907,32934,33016,33043,33233,33260,33342,33369,33451,33586,33668,33695,33777,33804,33885,33912,34103,34130,34211,34239,34320,34456,34537,34565,34646,34673,34755,34782,34972,34999,35081,35108,35190,35326,35407,35434,35516,35543,35624,35652,35842,35869,35951,35978,36059,36195,36277,36304,36385,36412,36494,36521,36711,36739,36820,36847,36929,37065,37146,37173,37255,37282,37364,37391,37581,37608,37690,37717,37798,37826,38016,38043,38124,38152,38233,38260,38451,38478,38559,38586,38668,38804,38885,38912,38994,39021,39103,39130,39320,39347,39429,39456,39537,39673,39755,39782,39864,39891,39972,39999,40190,40217,40298,40326,40407,40543,40624,40652,40733,40760,40842,40869,41059,41086,41168,41195,41277,41412,41494,41521,41603,41630,41711,41739,41929,41956,42037,42065,42146,42282,42364,42391,42472,42499,42581,42608,42798,42826,42907,42934,43016,43152,43233,43260,43342,43369,43451,43478,43668,43695,43777,43804,43885,44021,44103,44130,44211,44239,44320,44347,44537,44565,44646,44673,44755,44891,44972,44999,45081,45108,45190,45217,45407,45434,45516,45543,45624,45760,45842,45869,45951,45978,46059,46086,46277,46304,46385,46412,46494,46630,46711,46739,46820,46847,46929,46956,47146,47173,47255,47282,47364,47499,47581,47608,47690,47717,47798,47826,48016,48043,48124,48152,48233,48260,48451,48478,48559,48586,48668,48695,48885,48912,48994,49021,49103,49239,49320,49347,49429,49456,49537,49565,49755,49782,49864,49891,49972,50108,50190,50217,50298,50326,50407,50434,50624,50652,50733,50760,50842,50978,51059,51086,51168,51195,51277,51304,51494,51521,51603,51630,51711,51847,51929,51956,52037,52065,52146,52173,52364,52391,52472,52499,52581,52717,52798,52826,52907,52934,53016,53043,53233,53260,53342,53369,53451,53586,53668,53695,53777,53804,53885,53912,54103,54130,54211,54239,54320,54456,54537,54565,54646,54673,54755,54782,54972,54999,55081,55108,55190,55217,55407,55434,55516,55543,55624,55652,55842,55869,55951,55978,56059,56195,56277,56304,56385,56412,56494,56521,56711,56739,56820,56847,56929,57065,57146,57173,57255,57282,57364,57391,57581,57608,57690,57717,57798,57934,58016,58043,58124,58152,58233,58260,58451,58478,58559,58586,58668,58804,58885,58912,58994,59021,59103,59130,59320,59347,59429,59456,59537,59673,59755,59782,59864,59891,59972,59999,60190,60217,60298,60326,60407,60543,60624,60652,60733,60760,60842,60869,61059,61086,61168,61195,61277,61412,61494,61521,61603,61630,61711,61739,61929,61956,62037,62065,62146,62173,62364,62391,62472,62499,62581,62608,62798,62825,62907,62934,63016,63152,63233,63260,63342,63369,63450,63478,63668,63695,63777,63804,63885,64021,64103,64130,64211,64239,64320,64347,64537,64565,64646,64673,64755,64891,64972,64999,65081,65108,65190,65217,65407,65434,65516,65543,65624,65760,65842,65869,65950,65978,66059,66086,66277,66304,66385,66412,66494,66630,66711,66739,66820,66847,66929,66956,67146,67173,67255,67282,67364,67499,67581,67608,67690,67717,67798,67825,68016,68043,68124,68152,68233,68369,68450,68478,68559,68586,68668,68695,68885,68912,68994,69021,69103,69130,69320,69347,69429,69456,69537,69565,71277,71304,73016,73043,76494,76521,78233,78260,79972,79999,83450,83478,85190,85217,86929,86956,90407,90434,92146,92173,93885,93912,95624,96521,96929,96956,97363,97391,97581,97608,97690,97717,97798,97934,98016,98043,98124,98152,98233,98260,98450,98478,98559,98586,98668,98804,98885,98912,98994,99021,99103,99130,99320,99347,99429,99456,99537,99673,99755,99782,99863,99891,99972,99999,100190,100217,100298,100325,100407,100434,100624,100652,100733,100760,100842,100869,101059,101086,101168,101195,101277,101412,101494,101521,101603,101630,101711,101738,101929,101956,102037,102065,102146,102282,102363,102391,102472,102499,102581,102608,102798,102825,102907,102934,103016,103152,103233,103260,103342,103369,103450,103478,103668,103695,103777,103804,103885,103912,104103,104130,104211,104238,104320,104347,104537,104565,104646,104673,104755,104891,104972,104999,105081,105108,105190,105217,105407,105434,105516,105543,105624,105760,105842,105869,105950,105978,106059,106086,106277,106304,106385,106412,106494,106630,106711,106738,106820,106847,106929,106956,107146,107173,107255,107282,107363,107391,107581,107608,107690,107717,107798,107825,108016,108043,108124,108152,108233,108369,108450,108478,108559,108586,108668,108695,108885,108912,108994,109021,109103,109238,109320,109347,109429,109456,109537,109565,109755,109782,109863,109891,109972,110108,110190,110217,110298,110325,110407,110434,110570,110597,110733,110760,110842,110869,111005,111032,111168,111168,111277,111304,111494,111521,111603,111630,111711,111847,111929,111956,112037,112065,112146,112173,112363,112391,112472,112499,112581,112717,112798,112825,112907,112934,113016,113043,113233,113260,113342,113369,113450,113586,113668,113695,113777,113804,113885,113912,114103,114130,114211,114238,114320,114347,114537,114565,114646,114673,114755,114782,114972,114999,115081,115108,115190,115325,115407,115434,115516,115543,115624,115652,115842,115869,115950,115978,116059,116195,116277,116304,116385,116412,116494,116521,116711,116738,116820,116847,116929,117065,117146,117173,117255,117282,117363,117391,117581,117608,117690,117717,117798,117934,118016,118043,118124,118152,118233,118260,118450,118478,118559,118586,118668,118804,118885,118912,118994,119021,119103,119130,119320,119347,119429,119456,119537,119673,119755,119782,119863,119891,119972,119999,120190,120217,120298,120325,120407,120543,120624,120652,120733,120760,120842,120869,121059,121086,121168,121195,121277,121304,121494,121521,121603,121630,121711,121738,121929,121956,122037,122065,122146,122282,122363,122391,122472,122499,122581,122608,122798,122825,122907,122934,123016,123152,123233,123260,123342,123369,123450,123478,123668,123695,123777,123804,123885,124021,124103,124130,124211,124238,124320,124347,124537,124565,124646,124673,124755,124891,124972,124999,125081,125108,125190,125217,125407,125434,125516,125543,125624,125760,125842,125869,125950,125978,126059,126086,126276,126304,126385,126412,126494,126630,126711,126738,126820,126847,126929,126956,127146,127173,127255,127282,127363,127499,127581,127608,127690,127717,127798,127825,128016,128043,128124,128151,128233,128260,128450,128478,128559,128586,128668,128695,128885,128912,128994,129021,129103,129238,129320,129347,129429,129456,129537,129565,129755,129782,129863,129891,129972,130108,130190,130217,130298,130325,130407,130434,130624,130651,130733,130760,130842,130978,131059,131086,131168,131195,131276,131304,131494,131521,131603,131630,131711,131847,131929,131956,132037,132065,132146,132173,132363,132391,132472,132499,132581,132717,132798,132825,132907,132934,133016,133043,133233,133260,133342,133369,133450,133586,133668,133695,133776,133804,133885,133912,134103,134130,134211,134238,134320,134456,134537,134565,134646,134673,134755,134782,134972,134999,135081,135108,135190,135217,135407,135434,135516,135543,135624,135651,135842,135869,135950,135978,136059,136195,136276,136304,136385,136412,136494,136521,136711,136738,136820,136847,136929,137065,137146,137173,137255,137282,137363,137391,137581,137608,137690,137717,137798,137934,138016,138043,138124,138151,138233,138260,138450,138478,138559,138586,138668,138804,138885,138912,138994,139021,139103,139130,139320,139347,139429,139456,139537,139673,139755,139782,139863,139891,139972,139999,140190,140217,140298,140325,140407,140543,140624,140651,140733,140760,140842,140869,141059,141086,141168,141195,141276,141412,141494,141521,141603,141630,141711,141738,141929,141956,142037,142065,142146,142282,142363,142391,142472,142499,142581,142608,142798,142825,142907,142934,143016,143151,143233,143260,143342,143369,143450,143478,143668,143695,143776,143804,143885,144021,144103,144130,144211,144238,144320,144347,144537,144565,144646,144673,144755,144891,144972,144999,145081,145108,145190,145217,145407,145434,145516,145543,145624,145651,145842,145869,145950,145978,146059,146086,146276,146304,146385,146412,146494,146630,146711,146738,146820,146847,146929,146956,147146,147173,147255,147282,147363,147499,147581,147608,147690,147717,147798,147825,148016,148043,148124,148151,148233,148369,148450,148478,148559,148586,148668,148695,148885,148912,148994,149021,149103,149238,149320,149347,149429,149456,149537,149565,149755,149782,149863,149891,149972,150108,150190,150217,150298,150325,150407,150434,150624,150651,150733,150760,150842,150978,151059,151086,151168,151195,151276,151304,151494,151521,151603,151630,151711,151847,151929,151956,152037,152065,152146,152173,152363,152391,152472,152499,152581,152608,152798,152825,152907,152934,153016,153043,153233,153260,153342,153369,153450,153586,153668,153695,153776,153804,153885,153912,154103,154130,154211,154238,154320,154456,154537,154565,154646,154673,154755,154782,154972,154999,155081,155108,155189,155325,155407,155434,155516,155543,155624,155651,155842,155869,155950,155978,156059,156195,156276,156304,156385,156412,156494,156521,156711,156738,156820,156847,156929,157064,157146,157173,157255,157282,157363,157391,157581,157608,157689,157717,157798,157934,158016,158043,158124,158151,158233,158260,158450,158478,158559,158586,158668,158804,158885,158912,158994,159021,159103,159130,159320,159347,159429,159456,159537,159564,159755,159782,159863,159891,159972,159999,160189,160217,160298,160325,160407,160543,160624,160651,160733,160760,160842,160869,161059,161086,161168,161195,161276,161412,161494,161521,161603,161630,161711,161738,161929,161956,162037,162064,162146,162282,162363,162391,162472,162499,162581,162608,162798,162825,162907,162934,163016,163151,163233,163260,163342,163369,163450,163478,163668,163695,163776,163804,163885,164021,164103,164130,164211,164238,164320,164347,164537,164564,164646,164673,164755,164891,164972,164999,165081,165108,165189,165217,165407,165434,165516,165543,165624,165760,165842,165869,165950,165978,166059,166086,166276,166304,166385,166412,166494,166521,166711,166738,166820,166847,166929,166956,168668,168695,170407,170434,173885,173912,175624,175651,177363,177391,180842,180869,182581,182608,184320,184347,187798,187825,189537,189564,191276,191304,193016,199999,199999,200004
	};

	logic [31:0] m5[1880] = '{
		0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,30,0,34,0,38,0,30,0,34,0,38,0,30,0,34,0,38,0,30,0,34,0,38,0,51,0,46,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,77,0,92,0,51,0,92,0,103,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,36,0,36,0,73,0,73,0,58,0,73,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,30,0,30,0,61,0,61,0,58,0,61,0,30,0,30,0,61,0,61,0,58,0,61,0,34,0,34,0,69,0,69,0,61,0,69,0,34,0,34,0,69,0,69,0,61,0,69,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,38,0,38,0,77,0,77,0,69,0,77,0,51,0,92,0,103,0,46,0,77,0,92,0,32,0,36,0,41,0,32,0,36,0,41,0,32,0,36,0,41,0,32,0,36,0,41,0,0,0,0
	};

endmodule